**.subckt bgr_1 VDD VSS Vbgr_out
*.iopin VDD
*.iopin VSS
*.opin Vbgr_out
XM1 Vstartup Vbgr_out VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=40 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 Vstartup Vbgr_out VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 net8 Vp VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=80 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XQ1 VSS VSS net1 sky130_fd_pr__pnp_05v5_W3p40L3p40 m=24
XM4 net9 Vp VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=80 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XQ2 VSS VSS Vd1 sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
XM5 Vbgr_out Vp VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=80 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 Vp Vstartup net2 VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Vss VSS GND 0
Vdd VDD GND 3.3
XM7 net12 Vp VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=40 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 net4 Vd1 net3 VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=80 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM9 net3 net4 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM10 net13 net4 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=6 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2
XM11 net14 Vd1 net5 VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=80 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM12 net15 Vd2 net5 VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=80 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM13 net6 net6 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=40 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM14 Vp net6 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=4 W=40 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
Vc6 net7 VSS 0
.save  i(vc6)
Vc1 net8 Vd2 0
.save  i(vc1)
Vc2 net9 Vd1 0
.save  i(vc2)
Vc3 net10 VSS 0
.save  i(vc3)
Vc4 net11 VSS 0
.save  i(vc4)
Vc5 net12 net4 0
.save  i(vc5)
Vc7 net5 net13 0
.save  i(vc7)
Vc8 Vp net14 0
.save  i(vc8)
Vc9 net6 net15 0
.save  i(vc9)
Vc10 net2 Vd1 0
.save  i(vc10)
C1 VDD Vp 10p m=1
C2 Vbgr_out VSS 1p m=1
XR9 net11 Vd1 VSS sky130_fd_pr__res_xhigh_po W=0.35 L=16.72 mult=1 m=1
XR2 net10 Vd2 VSS sky130_fd_pr__res_xhigh_po W=0.35 L=16.72 mult=1 m=1
XR3 net1 Vd2 VSS sky130_fd_pr__res_xhigh_po W=0.35 L=2.562 mult=1 m=1
XR1 net7 Vbgr_out VSS sky130_fd_pr__res_xhigh_po W=0.35 L=13.6 mult=1 m=1
XM15 Vp Vstartup net16 VSS sky130_fd_pr__nfet_g5v0d10v5 L=1 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Vc11 net16 Vd2 0
.save  i(vc11)
**** begin user architecture code
** manual skywater pdks install (with patches applied)
* .lib /home/vaibhav/share/pdk/sky130A/libs.tech/ngspice/models/sky130.lib.spice tt

** opencircuitdesign pdks install
.lib /home/vaibhav/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /home/vaibhav/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

**** end user architecture code
**.ends
.GLOBAL VSS
.GLOBAL GND
.GLOBAL VDD
**** begin user architecture code


.option METHOD=GEAR CHGTOL=1e-15 TRTOL=1 RELTOL=0.0001 VNTOL=0.1u
.option savecurrents savevoltages
.control
save all
//set temp=125
//op
//dc temp -40 125 10
dc Vdd 0 3.3 0.01
//tran 100n 10u
save v(Vdd) v(vbgr_out)
plot v(vbgr_out) V(Vdd)
print v(Vbgr_out)
//save all
write  /home/vaibhav/sky130-example/bgr_1.raw
.endc


**** end user architecture code
.end
